library verilog;
use verilog.vl_types.all;
entity count is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        en              : in     vl_logic;
        clr             : in     vl_logic;
        data            : out    vl_logic_vector(3 downto 0);
        t               : out    vl_logic
    );
end count;
