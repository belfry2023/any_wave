library verilog;
use verilog.vl_types.all;
entity any_wave_vlg_tst is
end any_wave_vlg_tst;
